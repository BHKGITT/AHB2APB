class seqs extends uvm_sequence#(apb_xtn);

`uvm_object_utils(seqs)

function new(string name="seqs");
super.new(name);
endfunction

endclass

